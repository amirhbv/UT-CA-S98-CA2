`timescale 1ns / 1ns
module Inst_memory(
	input [9 :0] address,
	output[15:0] inst
);
	reg [15:0] mem[0:1023] ;
	initial begin
		for (integer i = 0 ; i < 1024 ; i = i + 1)
			mem[i] <= {4'b1110, 2'b01, 2'b01, 8'b01000000 } ;

		mem[0]  <= {4'b1110, 2'b01, 2'b01, 8'b00000000  }; 	// ANDI R1, R1, 0

		mem[1]  <= {4'b0000, 2'b00,       10'b0111110100}; 	// LOAD R0, 500
		mem[2]  <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[3]  <= {4'b0000, 2'b00,       10'b0111110101}; 	// LOAD R0, 501
		mem[4]  <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[5]  <= {4'b0000, 2'b00,       10'b0111110110}; 	// LOAD R0, 502
		mem[6]  <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[7]  <= {4'b0000, 2'b00,       10'b0111110111}; 	// LOAD R0, 503
		mem[8]  <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[9]  <= {4'b0000, 2'b00,       10'b0111111000}; 	// LOAD R0, 504
		mem[10] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[11] <= {4'b0000, 2'b00,       10'b0111111001}; 	// LOAD R0, 505
		mem[12] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[13] <= {4'b0000, 2'b00,       10'b0111111010}; 	// LOAD R0, 506
		mem[14] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[15] <= {4'b0000, 2'b00,       10'b0111111011}; 	// LOAD R0, 507
		mem[16] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[17] <= {4'b0000, 2'b00,       10'b0111111100}; 	// LOAD R0, 508
		mem[18] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[19] <= {4'b0000, 2'b00,       10'b0111111101}; 	// LOAD R0, 509
		mem[20] <= {4'b1000, 2'b01, 2'b00, 8'b00000010  }; 	// ADD  R1, R0

		mem[21] <= {4'b0001, 2'b01,       10'b0111111110}; 	// STORE R0, 510
	end

	assign inst = mem[address] ;
endmodule
